library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.kakeudon_fpu.all;

entity FDIV is
  Port (input1 : in  unsigned(31 downto 0);
        input2  : in  unsigned(31 downto 0);
        clk : in std_logic;
        output : out unsigned(31 downto 0));
end entity FDIV;

architecture RTL of FDIV is
  subtype unsigned_word is unsigned(31 downto 0);
  signal a, b: unsigned_word := (others => '0');
  signal a1, a2, a3, a4, a5: unsigned_word := (others => '0');
  signal inv_in, inv_out, ans: unsigned_word;
begin
  inv: FINV port map (
    input => b, clk => clk, output => inv_out
  );
  mul: FMUL_OLD port map (
    input1 => a5, input2 => inv_in, clk => clk, output => ans
  );
  a <= (others => 'X') when TO_01(input1, 'X')(0) = 'X' else
       input1(31)&(30 downto 0 => '0') when input1(30 downto 23) = x"00" else
       input1;
  b <= (others => 'X') when TO_01(input2, 'X')(0) = 'X' else
       input2(31)&(30 downto 0 => '0') when input2(30 downto 23) = x"00" else
       input2;
  output <= ans;

  fdiv_proc: process(input1, input2, clk)
  begin
    if rising_edge(clk) then
      a5 <= a4;
      a4 <= a3;
      a3 <= a2;
      a2 <= a1;
      a1 <= a;
      inv_in <= inv_out;
    end if;
  end process;
end architecture RTL;
